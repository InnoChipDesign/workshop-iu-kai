module multiplier # (
    parameter int DLEN = 3
) (
    input  [DLEN - 1:0] a,
    input  [DLEN - 1:0] b,

    output [DLEN - 1:0] out
);

endmodule
