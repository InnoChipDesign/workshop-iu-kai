module subtractor (
    input  [4:0] a,
    input  [4:0] b,

    output [5:0] out
);

endmodule
