module half_adder (
    input  a,
    input  b,

    output q,
    output carry_out
);

    // Task:
    // Implement a half adder module using basic logic gates (or, and, xor, not, etc.)

endmodule
