module equality (
    input  [4:0] a,
    input  [4:0] b,

    // output
);

endmodule
