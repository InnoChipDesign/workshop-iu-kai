module adder (
    input  a4, a3, a2, a1, a0,
    input  b4, b3, b2, b1, b0,

    output q5, q4, q3, q2, q1, q0
);

    // Task:
    // Implement 5-bit adder using half_adder and full_adder instances


endmodule
