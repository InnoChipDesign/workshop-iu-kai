module alu
(
    input  [4:0] a,
    input  [4:0] b,

    input  [1:0] opcode,

    output       overflow,
    output [4:0] result
);

endmodule
