module half_adder
(
    input  a,
    input  b,

    output q,
    output carry_out
);

    // Задание:
    // Реализовать модуль полусумматора используя логические элементы (or, and, xor, not, и т.д.)


endmodule
