module equality
(
    input  [4:0] a,
    input  [4:0] b,

    output       equal
);

    // Task:
    // Implement a 5-bit equality checker

endmodule
