module full_adder
(
    input  carry_in,
    input  a,
    input  b,

    output q,
    output carry_out
);

    // Task:
    // Implement a full adder module using half_adders

endmodule
