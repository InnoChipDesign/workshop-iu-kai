module adder
(
    input  a4, a3, a2, a1, a0,
    input  b4, b3, b2, b1, b0,

    output overflow,
    output q4, q3, q2, q1, q0
);

    // Задание:
    // Реализовать модуль 5-ти битного сумматора используя модули half_adder и full_adder


endmodule
