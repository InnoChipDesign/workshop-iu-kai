module subtractor
(
    input  [4:0] a,
    input  [4:0] b,

    output overflow,
    output [4:0] out
);

endmodule
