module full_adder
(
    input  carry_in,
    input  a,
    input  b,

    output q,
    output carry_out
);

    // Задание:
    // Реализовать модуль полного сумматора используя модули полусумматоров


endmodule
