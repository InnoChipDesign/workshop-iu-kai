module mux5bit
(
    input  [4:0] in0,
    input  [4:0] in1,
    input  [4:0] in2,
    input  [4:0] in3,

    input  [1:0] select,

    output [4:0] result
);

endmodule
